library IEEE;
use IEEE.STD_LOGIC_1164.all;

package constants is
    constant TEST: std_logic := '1';
end constants;