----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:28:24 11/17/2015 
-- Design Name: 
-- Module Name:    pc - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity pc is
    Port ( input : in  STD_LOGIC_VECTOR (15 downto 0);
           output : out  STD_LOGIC_VECTOR (15 downto 0);
           clk : in  STD_LOGIC;
           wr : in  STD_LOGIC;
			  rst : in STD_LOGIC);
end pc;

architecture Behavioral of pc is

begin
    process (clk, rst)
    begin
	     if (rst = '1') then
		      output <= (others=>'0');
		  elsif (falling_edge(clk))
        then
            if (wr = '1')
            then
                output <= input;
            end if;
         end if;
		
    end process;
end Behavioral;

